--****** FLIPFLOP SR****************************************************************


library ieee;
use ieee. std_logic_1164.all;
use ieee. std_logic_arith.all;
use ieee. std_logic_unsigned.all;
 
entity SR_FF is
PORT( 	S,R,CLOCK: in std_logic;
			Q: out std_logic);
end SR_FF;
 
Architecture behavioral of SR_FF is
begin
	PROCESS(CLOCK)
	variable tmp: std_logic;
	begin
		if(rising_edge(CLOCK)) then
			if(S='0' and R='0')then tmp:=tmp;
			elsif(S='1' and R='1')then tmp:='Z';
			elsif(S='0' and R='1')then tmp:='0';
			else tmp:='1';
			end if;
		end if;
		Q <= tmp;
	end PROCESS;
end behavioral;