library ieee;
use ieee.std_logic_1164.all;

entity practica2 is port(

);
end practica2;

architecture behavior of practica2 is
begin 



end behavior;
